
module cache #(
	parameter	WIDTH = 1
)(
	input logic 	clk,
	input logic 	rst
);

// Black box

endmodule